









module variableROM();

endmodule
